module test(in,clk,out)
input in,clk;
output out;
wire out;

assign out= 2*in;


endmodule
